-------------------------------------------------------------------------------
--                        VGA Controller - Project
-------------------------------------------------------------------------------
-- ENTITY:         io_logic
-- FILENAME:       io_logic_rtl_cfg.vhd
-- ARCHITECTURE:   rtl
-- ENGINEER:       Jonas Berger
-- DATE:           27.09.2022
-- VERSION:        1.0
-------------------------------------------------------------------------------
-- DESCRIPTION:    This is the configuration for the entity io_logic and the
--                 architecture rtl
-------------------------------------------------------------------------------
-- REFERENCES:     (none)
-------------------------------------------------------------------------------
-- PACKAGES:       (none)
-------------------------------------------------------------------------------
-- CHANGES:        Version 1.0 - JB - 27.09.2022
-------------------------------------------------------------------------------

configuration io_logic_rtl_cfg of io_logic is
    for rtl              -- architecture rtl is used for entity io_logic
    end for;
end io_logic_rtl_cfg;
