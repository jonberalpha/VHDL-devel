-------------------------------------------------------------------------------
--                        VGA Controller - Project
-------------------------------------------------------------------------------
-- ENTITY:         rom2_cntrl
-- FILENAME:       rom2_cntrl_rtl_cfg.vhd
-- ARCHITECTURE:   rtl
-- ENGINEER:       Jonas Berger
-- DATE:           01.10.2022
-- VERSION:        1.0
-------------------------------------------------------------------------------
-- DESCRIPTION:    This is the configuration for the entity rom2_cntrl and the
--                 architecture rtl
-------------------------------------------------------------------------------
-- REFERENCES:     (none)
-------------------------------------------------------------------------------
-- PACKAGES:       (none)
-------------------------------------------------------------------------------
-- CHANGES:        Version 1.0 - JB - 01.10.2022
-------------------------------------------------------------------------------

configuration rom2_cntrl_rtl_cfg of rom2_cntrl is
    for rtl              -- architecture rtl is used for entity rom2_cntrl
    end for;
end rom2_cntrl_rtl_cfg;
