configuration tb_mc8051_sim_cfg of tb_mc8051 is
  for sim
  end for;
end tb_mc8051_sim_cfg;
