-------------------------------------------------------------------------------
--                        Calculator - Project
-------------------------------------------------------------------------------
-- ENTITY:         calc_ctrl
-- FILENAME:       calc_ctrl_rtl_cfg.vhd
-- ARCHITECTURE:   rtl
-- ENGINEER:       Jonas Berger
-- DATE:           17.03.2022
-- VERSION:        1.0
-------------------------------------------------------------------------------
-- DESCRIPTION:    This is the configuration for the entity calc_ctrl and the
--                 architecture rtl.
-------------------------------------------------------------------------------
-- REFERENCES:     (none)
-------------------------------------------------------------------------------
-- PACKAGES:       (none)
-------------------------------------------------------------------------------
-- CHANGES:        Version 1.0 - JB - 17.03.2022
-------------------------------------------------------------------------------

configuration calc_ctrl_rtl_cfg of calc_ctrl is
  for rtl        -- architecture rtl is used for entity calc_ctrl
  end for;
end calc_ctrl_rtl_cfg;
