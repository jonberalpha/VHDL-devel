-------------------------------------------------------------------------------
--                        VGA Controller - Project
-------------------------------------------------------------------------------
-- ENTITY:         vga_cntrl
-- FILENAME:       vga_cntrl_rtl_cfg.vhd
-- ARCHITECTURE:   rtl
-- ENGINEER:       Jonas Berger
-- DATE:           19.03.2022
-- VERSION:        1.0
-------------------------------------------------------------------------------
-- DESCRIPTION:    This is the configuration for the entity vga_cntrl and the
--                 architecture rtl
-------------------------------------------------------------------------------
-- REFERENCES:     (none)
-------------------------------------------------------------------------------
-- PACKAGES:       (none)
-------------------------------------------------------------------------------
-- CHANGES:        Version 1.0 - JB - 19.09.2022
-------------------------------------------------------------------------------

configuration vga_cntrl_rtl_cfg of vga_cntrl is
    for rtl              -- architecture rtl is used for entity vga_cntrl
    end for;
end vga_cntrl_rtl_cfg;
