-------------------------------------------------------------------------------
--                        VGA Controller - Project
-------------------------------------------------------------------------------
-- ENTITY:         patgen1
-- FILENAME:       patgen1_rtl_cfg.vhd
-- ARCHITECTURE:   rtl
-- ENGINEER:       Jonas Berger
-- DATE:           28.09.2022
-- VERSION:        1.0
-------------------------------------------------------------------------------
-- DESCRIPTION:    This is the configuration for the entity patgen1 and the
--                 architecture rtl
-------------------------------------------------------------------------------
-- REFERENCES:     (none)
-------------------------------------------------------------------------------
-- PACKAGES:       (none)
-------------------------------------------------------------------------------
-- CHANGES:        Version 1.0 - JB - 28.09.2022
-------------------------------------------------------------------------------

configuration patgen1_rtl_cfg of patgen1 is
    for rtl              -- architecture rtl is used for entity patgen1
    end for;
end patgen1_rtl_cfg;
