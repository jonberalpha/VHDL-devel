-------------------------------------------------------------------------------
--                        VGA Controller - Project
-------------------------------------------------------------------------------
-- ENTITY:         src_mux
-- FILENAME:       src_mux_rtl_cfg.vhd
-- ARCHITECTURE:   rtl
-- ENGINEER:       Jonas Berger
-- DATE:           27.09.2022
-- VERSION:        1.0
-------------------------------------------------------------------------------
-- DESCRIPTION:    This is the configuration for the entity src_mux and the
--                 architecture rtl
-------------------------------------------------------------------------------
-- REFERENCES:     (none)
-------------------------------------------------------------------------------
-- PACKAGES:       (none)
-------------------------------------------------------------------------------
-- CHANGES:        Version 1.0 - JB - 27.09.2022
-------------------------------------------------------------------------------

configuration src_mux_rtl_cfg of src_mux is
    for rtl              -- architecture rtl is used for entity src_mux
    end for;
end src_mux_rtl_cfg;
