library ieee;
use ieee.std_logic_1164.all;

use std.textio.all;

entity tb_mc8051 is
end;
