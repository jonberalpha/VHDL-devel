-------------------------------------------------------------------------------
--                        VGA Controller - Project
-------------------------------------------------------------------------------
-- ENTITY:         rom1_cntrl
-- FILENAME:       rom1_cntrl_rtl_cfg.vhd
-- ARCHITECTURE:   rtl
-- ENGINEER:       Jonas Berger
-- DATE:           01.10.2022
-- VERSION:        1.0
-------------------------------------------------------------------------------
-- DESCRIPTION:    This is the configuration for the entity rom1_cntrl and the
--                 architecture rtl
-------------------------------------------------------------------------------
-- REFERENCES:     (none)
-------------------------------------------------------------------------------
-- PACKAGES:       (none)
-------------------------------------------------------------------------------
-- CHANGES:        Version 1.0 - JB - 01.10.2022
-------------------------------------------------------------------------------

configuration rom1_cntrl_rtl_cfg of rom1_cntrl is
    for rtl              -- architecture rtl is used for entity rom1_cntrl
    end for;
end rom1_cntrl_rtl_cfg;
